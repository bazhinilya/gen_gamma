module subtractor(a0, a1, a2, a3, a4, a5, a6, a7, a8, b0, b1, b2, b3,
     b4, b5, b6, b7, q0, q1, q2, q3, q4, q5, q6, q7);
  input a0, a1, a2, a3, a4, a5, a6, a7, a8, b0, b1, b2, b3, b4, b5, b6,
       b7;
  output q0, q1, q2, q3, q4, q5, q6, q7;
  wire a0, a1, a2, a3, a4, a5, a6, a7, a8, b0, b1, b2, b3, b4, b5, b6,
       b7;
  wire q0, q1, q2, q3, q4, q5, q6, q7;
  wire CARRY_IN, UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2,
       UNCONNECTED3, UNCONNECTED4, UNCONNECTED5;
  wire UNCONNECTED6, UNCONNECTED7, UNCONNECTED8, UNCONNECTED9,
       UNCONNECTED10, UNCONNECTED11, UNCONNECTED12, UNCONNECTED13;
  wire UNCONNECTED14, UNCONNECTED15, UNCONNECTED16, UNCONNECTED17,
       UNCONNECTED18, UNCONNECTED19, UNCONNECTED20, UNCONNECTED21;
  wire UNCONNECTED22, UNCONNECTED23, UNCONNECTED24, UNCONNECTED25,
       UNCONNECTED26, UNCONNECTED27, UNCONNECTED28, UNCONNECTED29;
  wire UNCONNECTED30, UNCONNECTED31, UNCONNECTED32, UNCONNECTED33,
       UNCONNECTED34, UNCONNECTED35, UNCONNECTED36, UNCONNECTED37;
  wire UNCONNECTED38, UNCONNECTED39, UNCONNECTED40, UNCONNECTED41,
       UNCONNECTED42, UNCONNECTED43, UNCONNECTED44, UNCONNECTED45;
  wire UNCONNECTED46, UNCONNECTED47, UNCONNECTED48, UNCONNECTED49,
       UNCONNECTED50, UNCONNECTED51, UNCONNECTED52, UNCONNECTED53;
  wire UNCONNECTED54, UNCONNECTED55, UNCONNECTED56, UNCONNECTED57,
       UNCONNECTED58, UNCONNECTED59, UNCONNECTED60, UNCONNECTED61;
  wire UNCONNECTED62, UNCONNECTED63, UNCONNECTED64, UNCONNECTED65,
       UNCONNECTED66, UNCONNECTED67, UNCONNECTED68, UNCONNECTED69;
  wire UNCONNECTED70, UNCONNECTED71, UNCONNECTED72, UNCONNECTED73,
       UNCONNECTED74, UNCONNECTED75, UNCONNECTED76, UNCONNECTED77;
  wire UNCONNECTED78, UNCONNECTED79, UNCONNECTED80, UNCONNECTED81,
       UNCONNECTED82, UNCONNECTED83, UNCONNECTED84, UNCONNECTED85;
  wire UNCONNECTED86, UNCONNECTED87, UNCONNECTED88, UNCONNECTED89,
       UNCONNECTED90, UNCONNECTED91, UNCONNECTED92, UNCONNECTED93;
  wire UNCONNECTED94, UNCONNECTED95, UNCONNECTED96, UNCONNECTED97,
       UNCONNECTED98, UNCONNECTED99, UNCONNECTED100, UNCONNECTED101;
  wire UNCONNECTED102, UNCONNECTED103, UNCONNECTED104, UNCONNECTED105,
       UNCONNECTED106, UNCONNECTED107, UNCONNECTED108, UNCONNECTED109;
  wire UNCONNECTED110, UNCONNECTED111, UNCONNECTED112, UNCONNECTED113,
       UNCONNECTED114, UNCONNECTED115, UNCONNECTED116, UNCONNECTED117;
  wire UNCONNECTED118, UNCONNECTED119, UNCONNECTED120, UNCONNECTED121,
       UNCONNECTED122, UNCONNECTED123, UNCONNECTED124, UNCONNECTED125;
  wire UNCONNECTED126, UNCONNECTED127, UNCONNECTED128, UNCONNECTED129,
       UNCONNECTED130, UNCONNECTED131, UNCONNECTED132, UNCONNECTED133;
  wire UNCONNECTED134, UNCONNECTED135, UNCONNECTED136, UNCONNECTED137,
       UNCONNECTED138, UNCONNECTED139, UNCONNECTED140, UNCONNECTED141;
  wire UNCONNECTED142, UNCONNECTED143, UNCONNECTED144, UNCONNECTED145,
       UNCONNECTED146, UNCONNECTED147, UNCONNECTED148, UNCONNECTED149;
  wire UNCONNECTED150, UNCONNECTED151, UNCONNECTED152, UNCONNECTED153,
       UNCONNECTED154, UNCONNECTED155, UNCONNECTED156, UNCONNECTED157;
  wire UNCONNECTED158, UNCONNECTED159, UNCONNECTED160, UNCONNECTED161,
       UNCONNECTED162, UNCONNECTED163, UNCONNECTED164, UNCONNECTED165;
  wire UNCONNECTED166, UNCONNECTED167, UNCONNECTED168, UNCONNECTED169,
       UNCONNECTED170, UNCONNECTED171, UNCONNECTED172, UNCONNECTED173;
  wire UNCONNECTED174, UNCONNECTED175, UNCONNECTED176, UNCONNECTED177,
       UNCONNECTED178, UNCONNECTED179, UNCONNECTED180, UNCONNECTED181;
  wire UNCONNECTED182, UNCONNECTED183, UNCONNECTED184, UNCONNECTED185,
       UNCONNECTED186, UNCONNECTED187, UNCONNECTED188, UNCONNECTED189;
  wire UNCONNECTED190, UNCONNECTED191, UNCONNECTED192, UNCONNECTED193,
       UNCONNECTED194, UNCONNECTED195, UNCONNECTED196, UNCONNECTED197;
  wire UNCONNECTED198, UNCONNECTED199, UNCONNECTED200, UNCONNECTED201,
       UNCONNECTED202, UNCONNECTED203, UNCONNECTED204, UNCONNECTED205;
  wire UNCONNECTED206, UNCONNECTED207, UNCONNECTED208, UNCONNECTED209,
       UNCONNECTED210, UNCONNECTED211, UNCONNECTED212, UNCONNECTED213;
  wire UNCONNECTED214, UNCONNECTED215, UNCONNECTED216, UNCONNECTED217,
       UNCONNECTED218, UNCONNECTED219, UNCONNECTED220, UNCONNECTED221;
  wire UNCONNECTED222, UNCONNECTED223, UNCONNECTED224, UNCONNECTED225,
       UNCONNECTED226, UNCONNECTED227, UNCONNECTED228, UNCONNECTED229;
  wire UNCONNECTED230, UNCONNECTED231, UNCONNECTED232, UNCONNECTED233,
       UNCONNECTED234, UNCONNECTED235, UNCONNECTED236, UNCONNECTED237;
  wire UNCONNECTED238, UNCONNECTED239, UNCONNECTED240, UNCONNECTED241,
       UNCONNECTED242, UNCONNECTED243, UNCONNECTED244, UNCONNECTED245;
  wire UNCONNECTED246, c1, c2, c3, c4, c5, c6, c7;
  wire g0, g1, g2, g3, g4, g5, g6, g7;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_16;
  wire n_17, n_18, n_19, n_20, n_21, p0, p1, p2;
  wire p3, p4, p5, p6, p7;
  assign CARRY_IN = 1'b1;
  full_sum dif0(.a (a0), .b ({UNCONNECTED29, UNCONNECTED28,
       UNCONNECTED27, UNCONNECTED26, UNCONNECTED25, UNCONNECTED24,
       UNCONNECTED23, UNCONNECTED22, UNCONNECTED21, UNCONNECTED20,
       UNCONNECTED19, UNCONNECTED18, UNCONNECTED17, UNCONNECTED16,
       UNCONNECTED15, UNCONNECTED14, UNCONNECTED13, UNCONNECTED12,
       UNCONNECTED11, UNCONNECTED10, UNCONNECTED9, UNCONNECTED8,
       UNCONNECTED7, UNCONNECTED6, UNCONNECTED5, UNCONNECTED4,
       UNCONNECTED3, UNCONNECTED2, UNCONNECTED1, UNCONNECTED0,
       UNCONNECTED, n_14}), .p0 (CARRY_IN), .q (q0), .g (g0), .p (p0));
  full_sum dif1(.a (a1), .b ({UNCONNECTED60, UNCONNECTED59,
       UNCONNECTED58, UNCONNECTED57, UNCONNECTED56, UNCONNECTED55,
       UNCONNECTED54, UNCONNECTED53, UNCONNECTED52, UNCONNECTED51,
       UNCONNECTED50, UNCONNECTED49, UNCONNECTED48, UNCONNECTED47,
       UNCONNECTED46, UNCONNECTED45, UNCONNECTED44, UNCONNECTED43,
       UNCONNECTED42, UNCONNECTED41, UNCONNECTED40, UNCONNECTED39,
       UNCONNECTED38, UNCONNECTED37, UNCONNECTED36, UNCONNECTED35,
       UNCONNECTED34, UNCONNECTED33, UNCONNECTED32, UNCONNECTED31,
       UNCONNECTED30, n_13}), .p0 (c1), .q (q1), .g (g1), .p (p1));
  full_sum dif2(.a (a2), .b ({UNCONNECTED91, UNCONNECTED90,
       UNCONNECTED89, UNCONNECTED88, UNCONNECTED87, UNCONNECTED86,
       UNCONNECTED85, UNCONNECTED84, UNCONNECTED83, UNCONNECTED82,
       UNCONNECTED81, UNCONNECTED80, UNCONNECTED79, UNCONNECTED78,
       UNCONNECTED77, UNCONNECTED76, UNCONNECTED75, UNCONNECTED74,
       UNCONNECTED73, UNCONNECTED72, UNCONNECTED71, UNCONNECTED70,
       UNCONNECTED69, UNCONNECTED68, UNCONNECTED67, UNCONNECTED66,
       UNCONNECTED65, UNCONNECTED64, UNCONNECTED63, UNCONNECTED62,
       UNCONNECTED61, n_10}), .p0 (c2), .q (q2), .g (g2), .p (p2));
  full_sum dif3(.a (a3), .b ({UNCONNECTED122, UNCONNECTED121,
       UNCONNECTED120, UNCONNECTED119, UNCONNECTED118, UNCONNECTED117,
       UNCONNECTED116, UNCONNECTED115, UNCONNECTED114, UNCONNECTED113,
       UNCONNECTED112, UNCONNECTED111, UNCONNECTED110, UNCONNECTED109,
       UNCONNECTED108, UNCONNECTED107, UNCONNECTED106, UNCONNECTED105,
       UNCONNECTED104, UNCONNECTED103, UNCONNECTED102, UNCONNECTED101,
       UNCONNECTED100, UNCONNECTED99, UNCONNECTED98, UNCONNECTED97,
       UNCONNECTED96, UNCONNECTED95, UNCONNECTED94, UNCONNECTED93,
       UNCONNECTED92, n_12}), .p0 (c3), .q (q3), .g (g3), .p (p3));
  full_sum dif4(.a (a4), .b ({UNCONNECTED153, UNCONNECTED152,
       UNCONNECTED151, UNCONNECTED150, UNCONNECTED149, UNCONNECTED148,
       UNCONNECTED147, UNCONNECTED146, UNCONNECTED145, UNCONNECTED144,
       UNCONNECTED143, UNCONNECTED142, UNCONNECTED141, UNCONNECTED140,
       UNCONNECTED139, UNCONNECTED138, UNCONNECTED137, UNCONNECTED136,
       UNCONNECTED135, UNCONNECTED134, UNCONNECTED133, UNCONNECTED132,
       UNCONNECTED131, UNCONNECTED130, UNCONNECTED129, UNCONNECTED128,
       UNCONNECTED127, UNCONNECTED126, UNCONNECTED125, UNCONNECTED124,
       UNCONNECTED123, n_11}), .p0 (c4), .q (q4), .g (g4), .p (p4));
  full_sum dif5(.a (a5), .b ({UNCONNECTED184, UNCONNECTED183,
       UNCONNECTED182, UNCONNECTED181, UNCONNECTED180, UNCONNECTED179,
       UNCONNECTED178, UNCONNECTED177, UNCONNECTED176, UNCONNECTED175,
       UNCONNECTED174, UNCONNECTED173, UNCONNECTED172, UNCONNECTED171,
       UNCONNECTED170, UNCONNECTED169, UNCONNECTED168, UNCONNECTED167,
       UNCONNECTED166, UNCONNECTED165, UNCONNECTED164, UNCONNECTED163,
       UNCONNECTED162, UNCONNECTED161, UNCONNECTED160, UNCONNECTED159,
       UNCONNECTED158, UNCONNECTED157, UNCONNECTED156, UNCONNECTED155,
       UNCONNECTED154, n_9}), .p0 (c5), .q (q5), .g (g5), .p (p5));
  full_sum dif6(.a (a6), .b ({UNCONNECTED215, UNCONNECTED214,
       UNCONNECTED213, UNCONNECTED212, UNCONNECTED211, UNCONNECTED210,
       UNCONNECTED209, UNCONNECTED208, UNCONNECTED207, UNCONNECTED206,
       UNCONNECTED205, UNCONNECTED204, UNCONNECTED203, UNCONNECTED202,
       UNCONNECTED201, UNCONNECTED200, UNCONNECTED199, UNCONNECTED198,
       UNCONNECTED197, UNCONNECTED196, UNCONNECTED195, UNCONNECTED194,
       UNCONNECTED193, UNCONNECTED192, UNCONNECTED191, UNCONNECTED190,
       UNCONNECTED189, UNCONNECTED188, UNCONNECTED187, UNCONNECTED186,
       UNCONNECTED185, n_8}), .p0 (c6), .q (q6), .g (g6), .p (p6));
  full_sum dif7(.a (a7), .b ({UNCONNECTED246, UNCONNECTED245,
       UNCONNECTED244, UNCONNECTED243, UNCONNECTED242, UNCONNECTED241,
       UNCONNECTED240, UNCONNECTED239, UNCONNECTED238, UNCONNECTED237,
       UNCONNECTED236, UNCONNECTED235, UNCONNECTED234, UNCONNECTED233,
       UNCONNECTED232, UNCONNECTED231, UNCONNECTED230, UNCONNECTED229,
       UNCONNECTED228, UNCONNECTED227, UNCONNECTED226, UNCONNECTED225,
       UNCONNECTED224, UNCONNECTED223, UNCONNECTED222, UNCONNECTED221,
       UNCONNECTED220, UNCONNECTED219, UNCONNECTED218, UNCONNECTED217,
       UNCONNECTED216, n_7}), .p0 (c7), .q (q7), .g (g7), .p (p7));
  INVXL g429(.A (b0), .Y (n_14));
  INVXL g428(.A (b1), .Y (n_13));
  INVXL g433(.A (b3), .Y (n_12));
  INVXL g431(.A (b4), .Y (n_11));
  INVXL g430(.A (b2), .Y (n_10));
  INVXL g432(.A (b5), .Y (n_9));
  INVXL g434(.A (b6), .Y (n_8));
  INVXL g435(.A (b7), .Y (n_7));
  XNOR2X1 g595__8780(.A (g6), .B (n_6), .Y (c7));
  NAND2XL g596__4296(.A (p6), .B (n_16), .Y (n_6));
  XNOR2X1 g597__3772(.A (g5), .B (n_5), .Y (n_16));
  NAND2XL g598__1474(.A (p5), .B (n_17), .Y (n_5));
  XNOR2X1 g599__4547(.A (g4), .B (n_4), .Y (n_17));
  NAND2XL g600__9682(.A (p4), .B (n_18), .Y (n_4));
  XNOR2X1 g601__2683(.A (g3), .B (n_3), .Y (n_18));
  NAND2XL g602__1309(.A (p3), .B (n_19), .Y (n_3));
  XNOR2X1 g603__6877(.A (g2), .B (n_2), .Y (n_19));
  NAND2XL g604__2900(.A (p2), .B (n_20), .Y (n_2));
  XNOR2X1 g605__2391(.A (g1), .B (n_1), .Y (n_20));
  NAND2XL g606__7675(.A (p1), .B (n_21), .Y (n_1));
  XNOR2X1 g607__7118(.A (g0), .B (n_0), .Y (n_21));
  NAND2XL g608__8757(.A (CARRY_IN), .B (p0), .Y (n_0));
  BUFX2 g609(.A (n_21), .Y (c1));
  BUFX2 g610(.A (n_20), .Y (c2));
  BUFX2 g611(.A (n_19), .Y (c3));
  BUFX2 g612(.A (n_18), .Y (c4));
  BUFX2 g613(.A (n_17), .Y (c5));
  BUFX2 g614(.A (n_16), .Y (c6));
endmodule

module gen_gamma_decoder(clk, rst_n, set0, set1, md, nk, od);
  input clk, rst_n, set0, set1;
  input [8:0] md;
  input [7:0] nk;
  output [7:0] od;
  wire clk, rst_n, set0, set1;
  wire [8:0] md;
  wire [7:0] nk;
  wire [7:0] od;
  wire [24:0] w;
  wire UNCONNECTED_HIER_Z;
  subtractor difference_two_list(.a0 (w[0]), .a1 (w[1]), .a2 (w[2]),
       .a3 (w[3]), .a4 (w[4]), .a5 (w[5]), .a6 (w[6]), .a7 (w[7]), .a8
       (UNCONNECTED_HIER_Z), .b0 (w[9]), .b1 (w[10]), .b2 (w[11]), .b3
       (w[12]), .b4 (w[13]), .b5 (w[14]), .b6 (w[15]), .b7 (w[16]), .q0
       (w[17]), .q1 (w[18]), .q2 (w[19]), .q3 (w[20]), .q4 (w[21]), .q5
       (w[22]), .q6 (w[23]), .q7 (w[24]));
  SDFFRHQX1 \saving_mix_data_q_reg[6] (.RN (rst_n), .CK (clk), .D
       (w[6]), .SI (md[6]), .SE (set0), .Q (w[6]));
  SDFFRHQX1 \saving_mix_data_q_reg[1] (.RN (rst_n), .CK (clk), .D
       (w[1]), .SI (md[1]), .SE (set0), .Q (w[1]));
  SDFFRHQX1 \saving_mix_data_q_reg[2] (.RN (rst_n), .CK (clk), .D
       (w[2]), .SI (md[2]), .SE (set0), .Q (w[2]));
  SDFFRHQX1 \saving_mix_data_q_reg[3] (.RN (rst_n), .CK (clk), .D
       (w[3]), .SI (md[3]), .SE (set0), .Q (w[3]));
  SDFFRHQX1 \saving_mix_data_q_reg[4] (.RN (rst_n), .CK (clk), .D
       (w[4]), .SI (md[4]), .SE (set0), .Q (w[4]));
  SDFFRHQX1 \saving_mix_data_q_reg[5] (.RN (rst_n), .CK (clk), .D
       (w[5]), .SI (md[5]), .SE (set0), .Q (w[5]));
  SDFFRHQX1 \saving_mix_data_q_reg[0] (.RN (rst_n), .CK (clk), .D
       (w[0]), .SI (md[0]), .SE (set0), .Q (w[0]));
  SDFFRHQX1 \saving_mix_data_q_reg[7] (.RN (rst_n), .CK (clk), .D
       (w[7]), .SI (md[7]), .SE (set0), .Q (w[7]));
  SDFFRHQX1 \saving_original_data_q_reg[3] (.RN (rst_n), .CK (clk), .D
       (od[3]), .SI (w[20]), .SE (set1), .Q (od[3]));
  SDFFRHQX1 \saving_original_data_q_reg[2] (.RN (rst_n), .CK (clk), .D
       (od[2]), .SI (w[19]), .SE (set1), .Q (od[2]));
  SDFFRHQX1 \saving_original_data_q_reg[1] (.RN (rst_n), .CK (clk), .D
       (od[1]), .SI (w[18]), .SE (set1), .Q (od[1]));
  SDFFRHQX1 \saving_original_data_q_reg[0] (.RN (rst_n), .CK (clk), .D
       (od[0]), .SI (w[17]), .SE (set1), .Q (od[0]));
  SDFFRHQX1 \saving_noise_key_q_reg[2] (.RN (rst_n), .CK (clk), .D
       (w[11]), .SI (nk[2]), .SE (set0), .Q (w[11]));
  SDFFRHQX1 \saving_original_data_q_reg[5] (.RN (rst_n), .CK (clk), .D
       (od[5]), .SI (w[22]), .SE (set1), .Q (od[5]));
  SDFFRHQX1 \saving_original_data_q_reg[6] (.RN (rst_n), .CK (clk), .D
       (od[6]), .SI (w[23]), .SE (set1), .Q (od[6]));
  SDFFRHQX1 \saving_original_data_q_reg[7] (.RN (rst_n), .CK (clk), .D
       (od[7]), .SI (w[24]), .SE (set1), .Q (od[7]));
  SDFFRHQX1 \saving_noise_key_q_reg[0] (.RN (rst_n), .CK (clk), .D
       (w[9]), .SI (nk[0]), .SE (set0), .Q (w[9]));
  SDFFRHQX1 \saving_noise_key_q_reg[1] (.RN (rst_n), .CK (clk), .D
       (w[10]), .SI (nk[1]), .SE (set0), .Q (w[10]));
  SDFFRHQX1 \saving_original_data_q_reg[4] (.RN (rst_n), .CK (clk), .D
       (od[4]), .SI (w[21]), .SE (set1), .Q (od[4]));
  SDFFRHQX1 \saving_noise_key_q_reg[3] (.RN (rst_n), .CK (clk), .D
       (w[12]), .SI (nk[3]), .SE (set0), .Q (w[12]));
  SDFFRHQX1 \saving_noise_key_q_reg[4] (.RN (rst_n), .CK (clk), .D
       (w[13]), .SI (nk[4]), .SE (set0), .Q (w[13]));
  SDFFRHQX1 \saving_noise_key_q_reg[5] (.RN (rst_n), .CK (clk), .D
       (w[14]), .SI (nk[5]), .SE (set0), .Q (w[14]));
  SDFFRHQX1 \saving_noise_key_q_reg[6] (.RN (rst_n), .CK (clk), .D
       (w[15]), .SI (nk[6]), .SE (set0), .Q (w[15]));
  SDFFRHQX1 \saving_noise_key_q_reg[7] (.RN (rst_n), .CK (clk), .D
       (w[16]), .SI (nk[7]), .SE (set0), .Q (w[16]));
endmodule

module top(clk_i, rst_n_i, set0_i, set1_i, md_i, nk_i, od_o);
  input clk_i, rst_n_i, set0_i, set1_i;
  input  [8:0] md_i;
  input  [7:0] nk_i;
  output [7:0] od_o;
  
  wire clk, rst_n, set0, set1;
  wire [7:0] od, nk;
  wire [8:0] md;
  
  wire VDDC, VDDO;
  wire VSSC, VSSO;
  
gen_gamma_decoder U1 (.clk(clk), 
  .rst_n(rst_n), 
  .set0(set0), 
  .set1(set1),  
  .md(md),
  .nk(nk), 
  .od(od)); 

PADDI PAD_clk   (.PAD(clk_i),   .Y(clk),   .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDI PAD_rst_n (.PAD(rst_n_i), .Y(rst_n), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDI PAD_set0  (.PAD(set0_i),  .Y(set0),  .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDI PAD_set1  (.PAD(set1_i),  .Y(set1),  .VDDIOR(VDDO), .VSSIOR(VSSO));

PADDO PAD_od0 (.PAD(od_o[0]), .A(od[0]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od1 (.PAD(od_o[1]), .A(od[1]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od2 (.PAD(od_o[2]), .A(od[2]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od3 (.PAD(od_o[3]), .A(od[3]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od4 (.PAD(od_o[4]), .A(od[4]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od5 (.PAD(od_o[5]), .A(od[5]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od6 (.PAD(od_o[6]), .A(od[6]), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADDO PAD_od7 (.PAD(od_o[7]), .A(od[7]), .VDDIOR(VDDO), .VSSIOR(VSSO));

PADDI PAD_md0 (.Y(md[0]), .PAD(md_i[0]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md1 (.Y(md[1]), .PAD(md_i[1]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md2 (.Y(md[2]), .PAD(md_i[2]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md3 (.Y(md[3]), .PAD(md_i[3]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md4 (.Y(md[4]), .PAD(md_i[4]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md5 (.Y(md[5]), .PAD(md_i[5]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md6 (.Y(md[6]), .PAD(md_i[6]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md7 (.Y(md[7]), .PAD(md_i[7]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_md8 (.Y(md[8]), .PAD(md_i[8]), .VDDIOR(VDDO), .VSSIOR(VSSO));

PADDI PAD_nk0 (.Y(nk[0]), .PAD(nk_i[0]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk1 (.Y(nk[1]), .PAD(nk_i[1]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk2 (.Y(nk[2]), .PAD(nk_i[2]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk3 (.Y(nk[3]), .PAD(nk_i[3]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk4 (.Y(nk[4]), .PAD(nk_i[4]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk5 (.Y(nk[5]), .PAD(nk_i[5]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk6 (.Y(nk[6]), .PAD(nk_i[6]), .VDDIOR(VDDO), .VSSIOR(VSSO)); 
PADDI PAD_nk7 (.Y(nk[7]), .PAD(nk_i[7]), .VDDIOR(VDDO), .VSSIOR(VSSO));

PADVDD PAD_VDD1 (.VDD(VDDC), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADVDD PAD_VDD2 (.VDD(VDDC), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADVDD PAD_VSS1 (.VSS(VSSC), .VDDIOR(VDDO), .VSSIOR(VSSO));
PADVDD PAD_VSS2 (.VSS(VSSC), .VDDIOR(VDDO), .VSSIOR(VSSO));

PADVDDIOR PAD_VDDIOR (.VDDIOR(VDDO), .VSSIOR(VSSO));
PADVSSIOR PAD_VSSIOR (.VDDIOR(VDDO), .VSSIOR(VSSO));

endmodule